LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.math_real.ceil;
USE ieee.math_real.log2;

PACKAGE general_package IS
    -- DATA FORMAT
    CONSTANT N_BITS : INTEGER := 8;
    CONSTANT N_FLOAT : INTEGER := 0;

    -- ARCHITECTURE PARAMETERS
    CONSTANT N_UNITS : INTEGER := 64; -- MUST BE A POWER OF TWO, SIZE OF THE NETWORK
    CONSTANT N_PARALL : INTEGER := 64; -- MUST BE A POWER OF TWO LESS THAN N_UNITS
    CONSTANT DEPTH : INTEGER := INTEGER(ceil(real(N_UNITS/N_PARALL)));

    -- ROM
    CONSTANT ADDRESS_WIDTH : INTEGER := INTEGER(ceil(log2(real(N_UNITS))));
    CONSTANT PARALL_WIDTH : INTEGER := INTEGER(ceil(log2(real(N_PARALL))));

    -- BUSES
    TYPE K_BUS IS ARRAY (N_PARALL - 1 DOWNTO 0) OF STD_LOGIC_VECTOR (N_BITS - 1 DOWNTO 0);
    TYPE N_BUS IS ARRAY (N_UNITS - 1 DOWNTO 0) OF STD_LOGIC_VECTOR (N_BITS - 1 DOWNTO 0);
    TYPE NK_BUS IS ARRAY (DEPTH - 1 DOWNTO 0) OF K_BUS;
END PACKAGE;